//
// LUT5 simulation model
//

module LUT5 #(
    parameter INIT_VALUE = "32'h00000000"
    ) (
    input A[4:0] ,
    output Y
  ) ;

//
// include user code here
//
  initial begin

  end

endmodule
