//
// LUT4 simulation model
//

module LUT4 #(
    parameter INIT_VALUE = "16'h0000"
    ) (
    input A[3:0] ,
    output Y
  ) ;

//
// include user code here
//
  initial begin

  end

endmodule
