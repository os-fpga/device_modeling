//
// CARRY_CHAIN simulation model
//

module CARRY_CHAIN (
    input P ,
    input G ,
    input CIN ,
    output O ,
    output COUT
  ) ;

//
// include user code here
//

endmodule
