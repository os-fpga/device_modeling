//
// LUT2 simulation model
//

module LUT2 #(
    parameter INIT_VALUE = "4'h0"
    ) (
    input A[1:0] ,
    output Y
  ) ;

//
// include user code here
//
  initial begin

  end

endmodule
