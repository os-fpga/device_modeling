//
// I_DDR simulation model
//

module I_DDR (
    input D ,
    input R ,
    input E ,
    input C ,
    output Q[1:0]
  ) ;

//
// include user code here
//

endmodule
