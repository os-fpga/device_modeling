//
// O_DDR simulation model
//

module O_DDR (
    input D[1:0] ,
    input R ,
    input E ,
    input C ,
    output Q
  ) ;

//
// include user code here
//

endmodule
