`timescale 1ns/1ps
`celldefine
//
// LATCHN simulation model
// Negative level-sensitive latch
//
// Copyright (c) 2023 Rapid Silicon, Inc.  All rights reserved.
//

module LATCHN (
  input D, // Data Input
  input G,
  output Q // Data Output
);

endmodule
`endcelldefine
