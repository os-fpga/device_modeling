//
// LUT6 simulation model
//

module LUT6 #(
    parameter INIT_VALUE = "64'h0000000000000000"
    ) (
    input A[5:0] ,
    output Y
  ) ;

//
// include user code here
//
  initial begin

  end

endmodule
