//
// O_DELAY simulation model
//

module O_DELAY #(
    parameter DELAY = "0"
    ) (
    input I ,
    input DLY_LOAD ,
    input DLY_ADJ ,
    input DLY_INCDEC ,
    output DLY_TAP_VALUE[5:0] ,
    output O
  ) ;

//
// include user code here
//
  initial begin

  end

endmodule
