//
// LUT1 simulation model
//

module LUT1 #(
    parameter INIT_VALUE = "2'h0"
    ) (
    input A ,
    output Y
  ) ;

//
// include user code here
//
  initial begin

  end

endmodule
