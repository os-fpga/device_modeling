`timescale 1ns/1ps
`celldefine
//
// LATCHR simulation model
// Positive level-sensitive latch with active-high asyncronous reset
//
// Copyright (c) 2023 Rapid Silicon, Inc.  All rights reserved.
//

module LATCHR (
  input D, // Data Input
  input G,
  input R, // Active-high asyncronous reset
  output Q // Data Output
);

endmodule
`endcelldefine
