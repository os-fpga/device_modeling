`timescale 1ns/1ps
`celldefine
//
// LATCH simulation model
// Positive level-sensitive latch
//
// Copyright (c) 2023 Rapid Silicon, Inc.  All rights reserved.
//

module LATCH (
  input D, // Data Input
  input G,
  output Q // Data Output
);

endmodule
`endcelldefine
