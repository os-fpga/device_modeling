//
// LUT3 simulation model
//

module LUT3 #(
    parameter INIT_VALUE = "8'h00"
    ) (
    input A[2:0] ,
    output Y
  ) ;

//
// include user code here
//
  initial begin

  end

endmodule
