//
// CLK_BUF simulation model
//

module CLK_BUF (
    input I ,
    output O
  ) ;

//
// include user code here
//

endmodule
